library ieee;
use ieee.std_logic_1164.all;

entity registrador is
port(clk, carga, reset : IN STD_LOGIC;
		   d : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		   q : OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END registrador;
ARCHITECTURE estrutura OF registrador IS
BEGIN
   PROCESS(clk, reset)
   BEGIN
      IF(reset = '1') THEN
          q <= "00000000";
      ELSIF(clk'EVENT AND clk = '1' AND carga = '1') THEN
          q <= d;
     END IF;
   END PROCESS;
END estrutura;

